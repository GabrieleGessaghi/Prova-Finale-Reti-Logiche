-- test prova 1
