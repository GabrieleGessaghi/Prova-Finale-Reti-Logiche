-- test prova 1
-- test prova 2